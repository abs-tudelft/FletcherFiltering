library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity FletcherWildcard is
  generic (
    BUS_ADDR_WIDTH : integer := 64
  );
  port (
    kcd_clk                     : in  std_logic;
    kcd_reset                   : in  std_logic;
    mmio_awvalid                : in  std_logic;
    mmio_awready                : out std_logic;
    mmio_awaddr                 : in  std_logic_vector(31 downto 0);
    mmio_wvalid                 : in  std_logic;
    mmio_wready                 : out std_logic;
    mmio_wdata                  : in  std_logic_vector(31 downto 0);
    mmio_wstrb                  : in  std_logic_vector(3 downto 0);
    mmio_bvalid                 : out std_logic;
    mmio_bready                 : in  std_logic;
    mmio_bresp                  : out std_logic_vector(1 downto 0);
    mmio_arvalid                : in  std_logic;
    mmio_arready                : out std_logic;
    mmio_araddr                 : in  std_logic_vector(31 downto 0);
    mmio_rvalid                 : out std_logic;
    mmio_rready                 : in  std_logic;
    mmio_rdata                  : out std_logic_vector(31 downto 0);
    mmio_rresp                  : out std_logic_vector(1 downto 0);
    ff_in_pkid_valid            : in  std_logic;
    ff_in_pkid_ready            : out std_logic;
    ff_in_pkid_dvalid           : in  std_logic;
    ff_in_pkid_last             : in  std_logic;
    ff_in_pkid                  : in  std_logic_vector(31 downto 0);
    ff_in_pkid_cmd_valid        : out std_logic;
    ff_in_pkid_cmd_ready        : in  std_logic;
    ff_in_pkid_cmd_firstIdx     : out std_logic_vector(31 downto 0);
    ff_in_pkid_cmd_lastidx      : out std_logic_vector(31 downto 0);
    ff_in_pkid_cmd_ctrl         : out std_logic_vector(bus_addr_width-1 downto 0);
    ff_in_pkid_cmd_tag          : out std_logic_vector(0 downto 0);
    ff_in_pkid_unl_valid        : in  std_logic;
    ff_in_pkid_unl_ready        : out std_logic;
    ff_in_pkid_unl_tag          : in  std_logic_vector(0 downto 0);
    ff_in_string1_valid         : in  std_logic;
    ff_in_string1_ready         : out std_logic;
    ff_in_string1_dvalid        : in  std_logic;
    ff_in_string1_last          : in  std_logic;
    ff_in_string1_length        : in  std_logic_vector(31 downto 0);
    ff_in_string1_count         : in  std_logic_vector(0 downto 0);
    ff_in_string1_chars_valid   : in  std_logic;
    ff_in_string1_chars_ready   : out std_logic;
    ff_in_string1_chars_dvalid  : in  std_logic;
    ff_in_string1_chars_last    : in  std_logic;
    ff_in_string1_chars_data    : in  std_logic_vector(7 downto 0);
    ff_in_string1_chars_count   : in  std_logic_vector(0 downto 0);
    ff_in_string1_cmd_valid     : out std_logic;
    ff_in_string1_cmd_ready     : in  std_logic;
    ff_in_string1_cmd_firstIdx  : out std_logic_vector(31 downto 0);
    ff_in_string1_cmd_lastidx   : out std_logic_vector(31 downto 0);
    ff_in_string1_cmd_ctrl      : out std_logic_vector(2*bus_addr_width-1 downto 0);
    ff_in_string1_cmd_tag       : out std_logic_vector(0 downto 0);
    ff_in_string1_unl_valid     : in  std_logic;
    ff_in_string1_unl_ready     : out std_logic;
    ff_in_string1_unl_tag       : in  std_logic_vector(0 downto 0);
    ff_in_string2_valid         : in  std_logic;
    ff_in_string2_ready         : out std_logic;
    ff_in_string2_dvalid        : in  std_logic;
    ff_in_string2_last          : in  std_logic;
    ff_in_string2_length        : in  std_logic_vector(31 downto 0);
    ff_in_string2_count         : in  std_logic_vector(0 downto 0);
    ff_in_string2_chars_valid   : in  std_logic;
    ff_in_string2_chars_ready   : out std_logic;
    ff_in_string2_chars_dvalid  : in  std_logic;
    ff_in_string2_chars_last    : in  std_logic;
    ff_in_string2_chars_data    : in  std_logic_vector(7 downto 0);
    ff_in_string2_chars_count   : in  std_logic_vector(0 downto 0);
    ff_in_string2_cmd_valid     : out std_logic;
    ff_in_string2_cmd_ready     : in  std_logic;
    ff_in_string2_cmd_firstIdx  : out std_logic_vector(31 downto 0);
    ff_in_string2_cmd_lastidx   : out std_logic_vector(31 downto 0);
    ff_in_string2_cmd_ctrl      : out std_logic_vector(2*bus_addr_width-1 downto 0);
    ff_in_string2_cmd_tag       : out std_logic_vector(0 downto 0);
    ff_in_string2_unl_valid     : in  std_logic;
    ff_in_string2_unl_ready     : out std_logic;
    ff_in_string2_unl_tag       : in  std_logic_vector(0 downto 0);
    ff_out_pkid_valid           : out std_logic;
    ff_out_pkid_ready           : in  std_logic;
    ff_out_pkid_dvalid          : out std_logic;
    ff_out_pkid_last            : out std_logic;
    ff_out_pkid                 : out std_logic_vector(31 downto 0);
    ff_out_pkid_cmd_valid       : out std_logic;
    ff_out_pkid_cmd_ready       : in  std_logic;
    ff_out_pkid_cmd_firstIdx    : out std_logic_vector(31 downto 0);
    ff_out_pkid_cmd_lastidx     : out std_logic_vector(31 downto 0);
    ff_out_pkid_cmd_ctrl        : out std_logic_vector(bus_addr_width-1 downto 0);
    ff_out_pkid_cmd_tag         : out std_logic_vector(0 downto 0);
    ff_out_pkid_unl_valid       : in  std_logic;
    ff_out_pkid_unl_ready       : out std_logic;
    ff_out_pkid_unl_tag         : in  std_logic_vector(0 downto 0);
    ff_out_string1_valid        : out std_logic;
    ff_out_string1_ready        : in  std_logic;
    ff_out_string1_dvalid       : out std_logic;
    ff_out_string1_last         : out std_logic;
    ff_out_string1_length       : out std_logic_vector(31 downto 0);
    ff_out_string1_count        : out std_logic_vector(0 downto 0);
    ff_out_string1_chars_valid  : out std_logic;
    ff_out_string1_chars_ready  : in  std_logic;
    ff_out_string1_chars_dvalid : out std_logic;
    ff_out_string1_chars_last   : out std_logic;
    ff_out_string1_chars_data   : out std_logic_vector(7 downto 0);
    ff_out_string1_chars_count  : out std_logic_vector(0 downto 0);
    ff_out_string1_cmd_valid    : out std_logic;
    ff_out_string1_cmd_ready    : in  std_logic;
    ff_out_string1_cmd_firstIdx : out std_logic_vector(31 downto 0);
    ff_out_string1_cmd_lastidx  : out std_logic_vector(31 downto 0);
    ff_out_string1_cmd_ctrl     : out std_logic_vector(2*bus_addr_width-1 downto 0);
    ff_out_string1_cmd_tag      : out std_logic_vector(0 downto 0);
    ff_out_string1_unl_valid    : in  std_logic;
    ff_out_string1_unl_ready    : out std_logic;
    ff_out_string1_unl_tag      : in  std_logic_vector(0 downto 0);
    ff_out_string2_valid        : out std_logic;
    ff_out_string2_ready        : in  std_logic;
    ff_out_string2_dvalid       : out std_logic;
    ff_out_string2_last         : out std_logic;
    ff_out_string2_length       : out std_logic_vector(31 downto 0);
    ff_out_string2_count        : out std_logic_vector(0 downto 0);
    ff_out_string2_chars_valid  : out std_logic;
    ff_out_string2_chars_ready  : in  std_logic;
    ff_out_string2_chars_dvalid : out std_logic;
    ff_out_string2_chars_last   : out std_logic;
    ff_out_string2_chars_data   : out std_logic_vector(7 downto 0);
    ff_out_string2_chars_count  : out std_logic_vector(0 downto 0);
    ff_out_string2_cmd_valid    : out std_logic;
    ff_out_string2_cmd_ready    : in  std_logic;
    ff_out_string2_cmd_firstIdx : out std_logic_vector(31 downto 0);
    ff_out_string2_cmd_lastidx  : out std_logic_vector(31 downto 0);
    ff_out_string2_cmd_ctrl     : out std_logic_vector(2*bus_addr_width-1 downto 0);
    ff_out_string2_cmd_tag      : out std_logic_vector(0 downto 0);
    ff_out_string2_unl_valid    : in  std_logic;
    ff_out_string2_unl_ready    : out std_logic;
    ff_out_string2_unl_tag      : in  std_logic_vector(0 downto 0)
  );
end entity;
architecture Implementation of FletcherWildcard is
begin
end architecture;
